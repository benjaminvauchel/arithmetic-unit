--*****************************************
--
-- Author: Benjamin
--
-- File: signed_nbit_adder_tb.vhd
--
-- Design units:
--	entity signed_nbit_adder_tb
--		function: check the acurracy of the nbit adder with signed type component
--	architecture tb_arch:
--		component: signed_nbit_adder
--			input: a_i, b_i
--			output: s_o
--		for statement implementation
--	configuration signed_nbit_adder_tb_conf
--		function: specify entity & architecture
--
-- Library
-- 	ieee.std_logic_1164: to use std_logic_vector, natural, boolean
--	LIB_RTL.design_pack
--
-- Synthesis and verification:
-- 	Synthesis software: ModelSim SE-64 10.6d
-- 	Options/Script:..
--	Target technology: ..
--
-- Revision history
--	version: 1.3
--	Date: 11/2023
--	Comments: Original
--
--******************************************

library IEEE;
use IEEE.std_logic_1164.all;

library lib_rtl;

entity signed_nbit_adder_tb is
    generic(nb_g : natural := 3);
end signed_nbit_adder_tb;

architecture tb_arch of signed_nbit_adder_tb is
  component signed_nbit_adder
    generic(nb_g : natural := nb_g);
    port(
      a_i, b_i : in std_logic_vector(nb_g-1 downto 0);
      s_o      : out std_logic_vector(nb_g downto 0));
end component;

  type sample is record
    a_i : std_logic_vector(nb_g-1 downto 0);
    b_i : std_logic_vector(nb_g-1 downto 0);
    s_o : std_logic_vector(nb_g downto 0);
  end record;
  type sample_array is array (natural range <>) of sample;

--  constant test_data: sample_array(255 downto 0) :=
--(("0000", "0000", "00000"), ("0000", "0001", "00001"), ("0000", "0010", "00010"), ("0000", "0011", "00011"), ("0000", "0100", "00100"), ("0000", "0101", "00101"), ("0000", "0110", "00110"), ("0000", "0111", "00111"), ("0000", "1000", "11000"), ("0000", "1001", "11001"), ("0000", "1010", "11010"), ("0000", "1011", "11011"), ("0000", "1100", "11100"), ("0000", "1101", "11101"), ("0000", "1110", "11110"), ("0000", "1111", "11111"), ("0001", "0000", "00001"), ("0001", "0001", "00010"), ("0001", "0010", "00011"), ("0001", "0011", "00100"), ("0001", "0100", "00101"), ("0001", "0101", "00110"), ("0001", "0110", "00111"), ("0001", "0111", "01000"), ("0001", "1000", "11001"), ("0001", "1001", "11010"), ("0001", "1010", "11011"), ("0001", "1011", "11100"), ("0001", "1100", "11101"), ("0001", "1101", "11110"), ("0001", "1110", "11111"), ("0001", "1111", "00000"), ("0010", "0000", "00010"), ("0010", "0001", "00011"), ("0010", "0010", "00100"), ("0010", "0011", "00101"), ("0010", "0100", "00110"), ("0010", "0101", "00111"), ("0010", "0110", "01000"), ("0010", "0111", "01001"), ("0010", "1000", "11010"), ("0010", "1001", "11011"), ("0010", "1010", "11100"), ("0010", "1011", "11101"), ("0010", "1100", "11110"), ("0010", "1101", "11111"), ("0010", "1110", "00000"), ("0010", "1111", "00001"), ("0011", "0000", "00011"), ("0011", "0001", "00100"), ("0011", "0010", "00101"), ("0011", "0011", "00110"), ("0011", "0100", "00111"), ("0011", "0101", "01000"), ("0011", "0110", "01001"), ("0011", "0111", "01010"), ("0011", "1000", "11011"), ("0011", "1001", "11100"), ("0011", "1010", "11101"), ("0011", "1011", "11110"), ("0011", "1100", "11111"), ("0011", "1101", "00000"), ("0011", "1110", "00001"), ("0011", "1111", "00010"), ("0100", "0000", "00100"), ("0100", "0001", "00101"), ("0100", "0010", "00110"), ("0100", "0011", "00111"), ("0100", "0100", "01000"), ("0100", "0101", "01001"), ("0100", "0110", "01010"), ("0100", "0111", "01011"), ("0100", "1000", "11100"), ("0100", "1001", "11101"), ("0100", "1010", "11110"), ("0100", "1011", "11111"), ("0100", "1100", "00000"), ("0100", "1101", "00001"), ("0100", "1110", "00010"), ("0100", "1111", "00011"), ("0101", "0000", "00101"), ("0101", "0001", "00110"), ("0101", "0010", "00111"), ("0101", "0011", "01000"), ("0101", "0100", "01001"), ("0101", "0101", "01010"), ("0101", "0110", "01011"), ("0101", "0111", "01100"), ("0101", "1000", "11101"), ("0101", "1001", "11110"), ("0101", "1010", "11111"), ("0101", "1011", "00000"), ("0101", "1100", "00001"), ("0101", "1101", "00010"), ("0101", "1110", "00011"), ("0101", "1111", "00100"), ("0110", "0000", "00110"), ("0110", "0001", "00111"), ("0110", "0010", "01000"), ("0110", "0011", "01001"), ("0110", "0100", "01010"), ("0110", "0101", "01011"), ("0110", "0110", "01100"), ("0110", "0111", "01101"), ("0110", "1000", "11110"), ("0110", "1001", "11111"), ("0110", "1010", "00000"), ("0110", "1011", "00001"), ("0110", "1100", "00010"), ("0110", "1101", "00011"), ("0110", "1110", "00100"), ("0110", "1111", "00101"), ("0111", "0000", "00111"), ("0111", "0001", "01000"), ("0111", "0010", "01001"), ("0111", "0011", "01010"), ("0111", "0100", "01011"), ("0111", "0101", "01100"), ("0111", "0110", "01101"), ("0111", "0111", "01110"), ("0111", "1000", "11111"), ("0111", "1001", "00000"), ("0111", "1010", "00001"), ("0111", "1011", "00010"), ("0111", "1100", "00011"), ("0111", "1101", "00100"), ("0111", "1110", "00101"), ("0111", "1111", "00110"), ("1000", "0000", "11000"), ("1000", "0001", "11001"), ("1000", "0010", "11010"), ("1000", "0011", "11011"), ("1000", "0100", "11100"), ("1000", "0101", "11101"), ("1000", "0110", "11110"), ("1000", "0111", "11111"), ("1000", "1000", "10000"), ("1000", "1001", "10001"), ("1000", "1010", "10010"), ("1000", "1011", "10011"), ("1000", "1100", "10100"), ("1000", "1101", "10101"), ("1000", "1110", "10110"), ("1000", "1111", "10111"), ("1001", "0000", "11001"), ("1001", "0001", "11010"), ("1001", "0010", "11011"), ("1001", "0011", "11100"), ("1001", "0100", "11101"), ("1001", "0101", "11110"), ("1001", "0110", "11111"), ("1001", "0111", "00000"), ("1001", "1000", "10001"), ("1001", "1001", "10010"), ("1001", "1010", "10011"), ("1001", "1011", "10100"), ("1001", "1100", "10101"), ("1001", "1101", "10110"), ("1001", "1110", "10111"), ("1001", "1111", "11000"), ("1010", "0000", "11010"), ("1010", "0001", "11011"), ("1010", "0010", "11100"), ("1010", "0011", "11101"), ("1010", "0100", "11110"), ("1010", "0101", "11111"), ("1010", "0110", "00000"), ("1010", "0111", "00001"), ("1010", "1000", "10010"), ("1010", "1001", "10011"), ("1010", "1010", "10100"), ("1010", "1011", "10101"), ("1010", "1100", "10110"), ("1010", "1101", "10111"), ("1010", "1110", "11000"), ("1010", "1111", "11001"), ("1011", "0000", "11011"), ("1011", "0001", "11100"), ("1011", "0010", "11101"), ("1011", "0011", "11110"), ("1011", "0100", "11111"), ("1011", "0101", "00000"), ("1011", "0110", "00001"), ("1011", "0111", "00010"), ("1011", "1000", "10011"), ("1011", "1001", "10100"), ("1011", "1010", "10101"), ("1011", "1011", "10110"), ("1011", "1100", "10111"), ("1011", "1101", "11000"), ("1011", "1110", "11001"), ("1011", "1111", "11010"), ("1100", "0000", "11100"), ("1100", "0001", "11101"), ("1100", "0010", "11110"), ("1100", "0011", "11111"), ("1100", "0100", "00000"), ("1100", "0101", "00001"), ("1100", "0110", "00010"), ("1100", "0111", "00011"), ("1100", "1000", "10100"), ("1100", "1001", "10101"), ("1100", "1010", "10110"), ("1100", "1011", "10111"), ("1100", "1100", "11000"), ("1100", "1101", "11001"), ("1100", "1110", "11010"), ("1100", "1111", "11011"), ("1101", "0000", "11101"), ("1101", "0001", "11110"), ("1101", "0010", "11111"), ("1101", "0011", "00000"), ("1101", "0100", "00001"), ("1101", "0101", "00010"), ("1101", "0110", "00011"), ("1101", "0111", "00100"), ("1101", "1000", "10101"), ("1101", "1001", "10110"), ("1101", "1010", "10111"), ("1101", "1011", "11000"), ("1101", "1100", "11001"), ("1101", "1101", "11010"), ("1101", "1110", "11011"), ("1101", "1111", "11100"), ("1110", "0000", "11110"), ("1110", "0001", "11111"), ("1110", "0010", "00000"), ("1110", "0011", "00001"), ("1110", "0100", "00010"), ("1110", "0101", "00011"), ("1110", "0110", "00100"), ("1110", "0111", "00101"), ("1110", "1000", "10110"), ("1110", "1001", "10111"), ("1110", "1010", "11000"), ("1110", "1011", "11001"), ("1110", "1100", "11010"), ("1110", "1101", "11011"), ("1110", "1110", "11100"), ("1110", "1111", "11101"), ("1111", "0000", "11111"), ("1111", "0001", "00000"), ("1111", "0010", "00001"), ("1111", "0011", "00010"), ("1111", "0100", "00011"), ("1111", "0101", "00100"), ("1111", "0110", "00101"), ("1111", "0111", "00110"), ("1111", "1000", "10111"), ("1111", "1001", "11000"), ("1111", "1010", "11001"), ("1111", "1011", "11010"), ("1111", "1100", "11011"), ("1111", "1101", "11100"), ("1111", "1110", "11101"), ("1111", "1111", "11110"));
constant test_data: sample_array(63 downto 0) := (
  ("000", "000", "0000"), ("000", "001", "0001"), ("000", "010", "0010"),
  ("000", "011", "0011"), ("000", "100", "1100"), ("000", "101", "1101"),
  ("000", "110", "1110"), ("000", "111", "1111"), ("001", "000", "0001"),
  ("001", "001", "0010"), ("001", "010", "0011"), ("001", "011", "0100"),
  ("001", "100", "1101"), ("001", "101", "1110"), ("001", "110", "1111"),
  ("001", "111", "0000"), ("010", "000", "0010"), ("010", "001", "0011"),
  ("010", "010", "0100"), ("010", "011", "0101"), ("010", "100", "1110"),
  ("010", "101", "1111"), ("010", "110", "0000"), ("010", "111", "0001"),
  ("011", "000", "0011"), ("011", "001", "0100"), ("011", "010", "0101"),
  ("011", "011", "0110"), ("011", "100", "1111"), ("011", "101", "0000"),
  ("011", "110", "0001"), ("011", "111", "0010"), ("100", "000", "1100"),
  ("100", "001", "1101"), ("100", "010", "1110"), ("100", "011", "1111"),
  ("100", "100", "1000"), ("100", "101", "1001"), ("100", "110", "1010"),
  ("100", "111", "1011"), ("101", "000", "1101"), ("101", "001", "1110"),
  ("101", "010", "1111"), ("101", "011", "0000"), ("101", "100", "1001"),
  ("101", "101", "1010"), ("101", "110", "1011"), ("101", "111", "1100"),
  ("110", "000", "1110"), ("110", "001", "1111"), ("110", "010", "0000"),
  ("110", "011", "0001"), ("110", "100", "1010"), ("110", "101", "1011"),
  ("110", "110", "1100"), ("110", "111", "1101"), ("111", "000", "1111"),
  ("111", "001", "0000"), ("111", "010", "0001"), ("111", "011", "0010"),
  ("111", "100", "1011"), ("111", "101", "1100"), ("111", "110", "1101"),
  ("111", "111", "1110")
);

	signal a_s, b_s: std_logic_vector(nb_g-1 downto 0);
  signal s_s: std_logic_vector(nb_g downto 0);
  signal test_ok: boolean := true;

begin

  process
    begin
      for i in test_data'range loop
        a_s <= test_data(i).a_i;
        b_s <= test_data(i).b_i;
        wait for 10 ns;

        if (s_s /= test_data(i).s_o) then
          test_ok <= false;
        else
          test_ok <= true;
        end if;

        assert (s_s = test_data(i).s_o)
        report "OUTPUT s_o WRONG."
        severity error;
        
      end  loop;
    wait;
  end process;

  DUT: signed_nbit_adder port map(a_s, b_s, s_s);

end architecture tb_arch;


configuration signed_nbit_adder_tb_conf of signed_nbit_adder_tb is
  for tb_arch
    for all: signed_nbit_adder
      use entity lib_rtl.signed_nbit_adder(struct_arch);
    end for;
  end for;
end configuration signed_nbit_adder_tb_conf;
